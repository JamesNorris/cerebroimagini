module dsp_main_tb;

endmodule